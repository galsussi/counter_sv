class transaction;
rand bit enable, load;
rand bit [7:0] Data_in ;
bit [7:0] count;
    function void display(string name);
    $display ("-----------------------------------------------------------");
    $display ("-%s-", name);
    $display ("-----------------------------------------------------------");
    $display ("-enable = %d , -load =%d ,-Data_in = %d", enable, load, Data_in);
    $display ("-count =%d", count);
    $display ("-----------------------------------------------------------");
            
    endfunction
endclass